Resistor bridge

.OP
VIN      1  0 10
L1       1  0 5n
R1       1  2 2
R2       1  3 1
R3       2  0 1
R4       3  0 2
R5       3  2 2
.END