Resistor bridge

.OP
VIN      1  0 10
R1       1  21 2
V1       21 2 0
R2       1  3 1
V3       2  22  0
R3       22  0 1
R4       3  0 2
R5       3  23 2
V5       23 2 0
.END
