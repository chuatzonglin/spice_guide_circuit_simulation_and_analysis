Resistor bridge

.OP
VIN      1  0 10
R1       1  21 2
V1       21 2 0
R2       1  31 1
V2       31 3 0
R3       22  0 1
V3       2  22  0
R4       33  30 2
C4       30  0  30p
V4       33 3 0
R5       3  23 2
V5       23 2 0
.END
