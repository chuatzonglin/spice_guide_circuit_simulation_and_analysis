Resistor divider
VIN	1	0	2volt
R1	1	2	4ohm
R2	2	0	1ohm
.SENS V(2)
.END
