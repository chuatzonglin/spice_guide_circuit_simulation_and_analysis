Resistor Bridge
Vin	1	0	1
R1	1	2	10
R2	1	3	2
R3	2	0	1
R4	3	0	5
R5	2	3	0.6
.DC	Vin 1	2	.1
.PRINT DC V(R1)
.PRINT DC V(2,3) V(3,2)
.PRINT DC I(R1)
.END